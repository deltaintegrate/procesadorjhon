----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:47:28 04/19/2018 
-- Design Name: 
-- Module Name:    mulx - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mulx is
    Port ( Amux : in  STD_LOGIC_VECTOR (31 downto 0);
           Bmux : in  STD_LOGIC_VECTOR (31 downto 0);
           sel : in  STD_LOGIC;
           Omux : out  STD_LOGIC_VECTOR (31 downto 0));
end mulx;

architecture Behavioral of mulx is

begin

	Omux <= Amux when (sel = '1') else Bmux;


end Behavioral;

